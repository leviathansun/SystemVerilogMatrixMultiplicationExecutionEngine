module ExecEngine (dataOut, dataInBus, clk, multRW, tranRW, memRW, subRW, addRW, multFleg, tranFleg, memFleg, subFleg, addFleg);
output reg [255:0] dataOut;
output reg fleg;

input [255:0] dataInBus;

always @ (posedge clk)
	


endmodule
module ExecEngine (dataOut, dataInBus, fleg);

endmodule
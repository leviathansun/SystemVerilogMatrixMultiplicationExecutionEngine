module ExecEngine (dataOut, dataInBus, fleg);
output reg [255:0] dataOut;
output reg fleg;

input [255:0] dataInBus;




endmodule